
-- Translatiing the VELO scrambler into VHDL from Verilog
-- Author Ben Jeffrey
-- Date Created 29/10/15
-- Algorithm by Sandeep from NIKHEF


-- IEEE VHDL standard library:
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VeloPixScrambler is
  port(
    dataIn      : in std_logic_vector(29 downto 0);
    state       : in std_logic_vector(29 downto 0);
    nextState   : out std_logic_vector(29 downto 0);
    dataOutEval : out std_logic_vector(29 downto 0)
    );
end VeloPixScrambler;

architecture a of VeloPixScrambler is

  signal myState : std_logic_vector(29 downto 0);
  
-------------------ALGORITHM ---------------------
begin

  myState(0)  <= dataIn(0)  XOR state(0)  XOR state(1)  XOR state(15)    XOR state(16);
  myState(1)  <= dataIn(1)  XOR state(1)  XOR state(2)  XOR state(16)    XOR state(17);
  myState(2)  <= dataIn(2)  XOR state(2)  XOR state(3)  XOR state(17)    XOR state(18);
  myState(3)  <= dataIn(3)  XOR state(3)  XOR state(4)  XOR state(18)    XOR state(19);
  myState(4)  <= dataIn(4)  XOR state(4)  XOR state(5)  XOR state(19)    XOR state(20);
  myState(5)  <= dataIn(5)  XOR state(5)  XOR state(6)  XOR state(20)    XOR state(21);
  myState(6)  <= dataIn(6)  XOR state(6)  XOR state(7)  XOR state(21)    XOR state(22);
  myState(7)  <= dataIn(7)  XOR state(7)  XOR state(8)  XOR state(22)    XOR state(23);
  myState(8)  <= dataIn(8)  XOR state(8)  XOR state(9)  XOR state(23)    XOR state(24);
  myState(9)  <= dataIn(9)  XOR state(9)  XOR state(10) XOR state(24)    XOR state(25);
  myState(10) <= dataIn(10) XOR state(10) XOR state(11) XOR state(25)    XOR state(26);
  myState(11) <= dataIn(11) XOR state(11) XOR state(12) XOR state(26)    XOR state(27);
  myState(12) <= dataIn(12) XOR state(12) XOR state(13) XOR state(27)    XOR state(28);
  myState(13) <= dataIn(13) XOR state(13) XOR state(14) XOR state(28)    XOR state(29);
  myState(14) <= dataIn(14) XOR state(14) XOR state(15) XOR state(29)    XOR myState(0);
  myState(15) <= dataIn(15) XOR state(15) XOR state(16) XOR myState(0) XOR myState(1);
  myState(16) <= dataIn(16) XOR state(16) XOR state(17) XOR myState(1) XOR myState(2);
  myState(17) <= dataIn(17) XOR state(17) XOR state(18) XOR myState(2) XOR myState(3);
  myState(18) <= dataIn(18) XOR state(18) XOR state(19) XOR myState(3) XOR myState(4);
  myState(19) <= dataIn(19) XOR state(19) XOR state(20) XOR myState(4) XOR myState(5);
  myState(20) <= dataIn(20) XOR state(20) XOR state(21) XOR myState(5) XOR myState(6);
  myState(21) <= dataIn(21) XOR state(21) XOR state(22) XOR myState(6) XOR myState(7);
  myState(22) <= dataIn(22) XOR state(22) XOR state(23) XOR myState(7) XOR myState(8);
  myState(23) <= dataIn(23) XOR state(23) XOR state(24) XOR myState(8) XOR myState(9);
  myState(24) <= dataIn(24) XOR state(24) XOR state(25) XOR myState(9) XOR myState(10);
  myState(25) <= dataIn(25) XOR state(25) XOR state(26) XOR myState(10) XOR myState(11);
  myState(26) <= dataIn(26) XOR state(26) XOR state(27) XOR myState(11) XOR myState(12);
  myState(27) <= dataIn(27) XOR state(27) XOR state(28) XOR myState(12) XOR myState(13);
  myState(28) <= dataIn(28) XOR state(28) XOR state(29) XOR myState(13) XOR myState(14);
  myState(29) <= dataIn(29) XOR state(29) XOR myState(0) XOR myState(14) XOR myState(15);

  dataOutEval <= myState;	
  nextState <= myState;

end a;
